/****************************************************************************
 * seq_item.svh
 ****************************************************************************/

/**
 * Class: seq_item
 * 
 * TODO: Add class documentation
 */
class seq_item extends uvm_object;
	`uvm_object_utils(seq_item)

	rand bit[7:0]		a;
	rand bit[7:0]		b;
	rand bit[7:0]		c;


endclass



