/****************************************************************************
 * uvm_rand_factory_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: uvm_rand_factory_pkg
 * 
 * TODO: Add package documentation
 */
package uvm_rand_factory_pkg;
	import uvm_pkg::*;

	`include "uvm_randomizer.svh"
	`include "uvm_randomizer_factory.svh"
	
	`include "uvm_rand_factory.svh"
`include "infact_uvm_randomizer_base.svh"
endpackage


