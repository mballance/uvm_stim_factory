

`include "uvm_macros.svh"
package uvm_stim_factory_tests_pkg;
	import uvm_pkg::*;
	import uvm_stim_factory_env_pkg::*;
	import uvm_stim_factory_pkg::*;

	`include "test_seq_item.svh"
	`include "test_seq_item2.svh"
	`include "test_seq_item_gen1.svh"
	`include "uvm_stim_factory_test_base.svh"
	`include "uvm_stim_factory_simple_override_test.svh"
	
endpackage
