
`include "uvm_macros.svh"

package uvm_stim_factory_env_pkg;
	import uvm_pkg::*;

	`include "uvm_stim_factory_env.svh"
	
endpackage
