/****************************************************************************
 * test_seq_item.svh
 ****************************************************************************/

/**
 * Class: test_seq_item
 * 
 * TODO: Add class documentation
 */
class test_seq_item extends uvm_sequence_item;
	`uvm_object_utils(test_seq_item)

	rand bit[3:0]	a, b, c;

endclass


