/****************************************************************************
 * seq_item_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: seq_item_pkg
 * 
 * TODO: Add package documentation
 */
package seq_item_pkg;
	import uvm_pkg::*;
	
	`include "seq_item.svh"

endpackage


