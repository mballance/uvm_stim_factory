/****************************************************************************
 * uvm_stim_factory_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"

/**
 * Package: uvm_stim_factory_pkg
 * 
 * TODO: Add package documentation
 */
package uvm_stim_factory_pkg;
	import uvm_pkg::*;

	`include "uvm_stim_gen.svh"
	`include "uvm_stim_factory.svh"
	`include "uvm_stim.svh"

endpackage


