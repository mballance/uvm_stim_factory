/****************************************************************************
 * uvm_stim_factory_tb.sv
 ****************************************************************************/

/**
 * Module: uvm_stim_factory_tb
 * 
 * TODO: Add module documentation
 */
`include "uvm_macros.svh"
module uvm_stim_factory_tb;
	import uvm_pkg::*;
	import uvm_stim_factory_tests_pkg::*;
	
	initial begin
		run_test();
	end

endmodule

