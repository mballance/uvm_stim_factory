/****************************************************************************
 * test_seq_item.svh
 ****************************************************************************/

/**
 * Class: test_seq_item
 * 
 * TODO: Add class documentation
 */
class test_seq_item2 extends test_seq_item;
	`uvm_object_utils(test_seq_item2)

endclass


