/****************************************************************************
 * seq_item_gen_pkg.sv
 ****************************************************************************/
`include "uvm_macros.svh"
`include "uvm_stim_macros.svh"

/**
 * Package: seq_item_gen_pkg
 * 
 * TODO: Add package documentation
 */
package seq_item_gen_pkg;
	import uvm_pkg::*;
	import seq_item_pkg::*;
	import uvm_stim_factory_pkg::*;

	`include "seq_item_gen.svh"

endpackage


